* SPICE3 file created from xor_2.ext - technology: scmos

.include "0.25-models"
.option scale=1u

M1000 out b a_16_31# Vdd CMOSP w=20 l=2
+  ad=240 pd=104 as=120 ps=52
M1001 a_n8_n28# b gnd gnd CMOSN w=8 l=2
+  ad=144 pd=84 as=96 ps=68
M1002 a_0_31# a out Vdd CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1003 a_n56_n48# b gnd gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1004 Vdd a_n56_n48# a_0_31# Vdd CMOSP w=20 l=2
+  ad=240 pd=116 as=0 ps=0
M1005 a_16_31# a_n25_n25# Vdd Vdd CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 out a a_n8_n28# gnd CMOSN w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1007 gnd a_n25_n25# a_n8_n28# gnd CMOSN w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_n25_n25# a Vdd Vdd CMOSP w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1009 a_n8_n28# a_n56_n48# out gnd CMOSN w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 a_n56_n48# b Vdd Vdd CMOSP w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1011 a_n25_n25# a gnd gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
C0 gnd a_n25_n25# 6.09fF
C1 Vdd b 4.77fF
C2 a_n8_n28# gnd 4.89fF
C3 gnd a_n56_n48# 21.73fF
C4 Vdd a_n25_n25# 12.20fF
C5 gnd a 7.15fF
C6 Vdd a_n56_n48# 3.76fF
C7 Vdd a 13.22fF
C8 Vdd out 5.88fF
C9 gnd b 12.62fF
C10 a_n8_n28# 0 2.82fF
C11 out 0 13.11fF
C12 b 0 30.07fF
C13 a_n25_n25# 0 16.61fF
C14 a_n56_n48# 0 16.61fF
C15 a 0 23.42fF
