magic
tech scmos
timestamp 1671730514
<< pwell >>
rect -75 -49 49 -19
rect -74 -59 49 -49
rect -75 -64 49 -59
rect -75 -69 47 -64
<< nwell >>
rect -75 20 49 65
<< polysilicon >>
rect -2 51 0 53
rect 6 51 8 53
rect 14 51 16 53
rect 22 51 24 53
rect -24 49 -22 51
rect -58 31 -56 33
rect -58 -44 -56 21
rect -24 -21 -22 39
rect -2 -20 0 31
rect 6 -20 8 31
rect 14 17 16 31
rect 14 -20 16 12
rect 22 1 24 31
rect 22 -20 24 -3
rect -24 -27 -22 -25
rect -58 -60 -56 -48
rect -2 -61 0 -28
rect 6 -39 8 -28
rect 6 -61 8 -43
rect 14 -61 16 -28
rect 22 -61 24 -28
<< ndiffusion >>
rect -8 -21 -2 -20
rect -30 -25 -29 -21
rect -25 -25 -24 -21
rect -22 -25 -21 -21
rect -17 -25 -16 -21
rect -8 -27 -7 -21
rect -3 -27 -2 -21
rect -8 -28 -2 -27
rect 0 -21 6 -20
rect 0 -27 1 -21
rect 5 -27 6 -21
rect 0 -28 6 -27
rect 8 -21 14 -20
rect 8 -27 9 -21
rect 13 -27 14 -21
rect 8 -28 14 -27
rect 16 -21 22 -20
rect 16 -27 17 -21
rect 21 -27 22 -21
rect 16 -28 22 -27
rect 24 -21 30 -20
rect 24 -27 25 -21
rect 29 -27 30 -21
rect 24 -28 30 -27
rect -64 -48 -63 -44
rect -59 -48 -58 -44
rect -56 -48 -55 -44
rect -51 -48 -49 -44
<< pdiffusion >>
rect -8 50 -2 51
rect -30 48 -24 49
rect -30 40 -29 48
rect -25 40 -24 48
rect -30 39 -24 40
rect -22 48 -16 49
rect -22 40 -21 48
rect -17 40 -16 48
rect -22 39 -16 40
rect -8 46 -7 50
rect -3 46 -2 50
rect -8 43 -2 46
rect -8 39 -7 43
rect -3 39 -2 43
rect -64 30 -58 31
rect -64 22 -63 30
rect -59 22 -58 30
rect -64 21 -58 22
rect -56 30 -50 31
rect -56 22 -55 30
rect -51 22 -50 30
rect -56 21 -50 22
rect -8 36 -2 39
rect -8 32 -7 36
rect -3 32 -2 36
rect -8 31 -2 32
rect 0 50 6 51
rect 0 46 1 50
rect 5 46 6 50
rect 0 43 6 46
rect 0 39 1 43
rect 5 39 6 43
rect 0 36 6 39
rect 0 32 1 36
rect 5 32 6 36
rect 0 31 6 32
rect 8 50 14 51
rect 8 46 9 50
rect 13 46 14 50
rect 8 43 14 46
rect 8 39 9 43
rect 13 39 14 43
rect 8 36 14 39
rect 8 32 9 36
rect 13 32 14 36
rect 8 31 14 32
rect 16 50 22 51
rect 16 46 17 50
rect 21 46 22 50
rect 16 43 22 46
rect 16 39 17 43
rect 21 39 22 43
rect 16 36 22 39
rect 16 32 17 36
rect 21 32 22 36
rect 16 31 22 32
rect 24 50 30 51
rect 24 46 25 50
rect 29 46 30 50
rect 24 43 30 46
rect 24 39 25 43
rect 29 39 30 43
rect 24 36 30 39
rect 24 32 25 36
rect 29 32 30 36
rect 24 31 30 32
<< metal1 >>
rect -67 58 -63 62
rect -59 58 37 62
rect 41 58 45 62
rect -63 30 -59 58
rect -29 48 -25 58
rect 9 50 13 58
rect -42 26 -38 30
rect -34 26 -28 30
rect -75 -1 -71 3
rect -67 -1 -62 3
rect -55 -39 -51 22
rect -43 12 -30 17
rect -21 -5 -17 40
rect -7 43 -3 46
rect 9 43 13 46
rect 25 43 29 46
rect -7 36 -3 39
rect 9 36 13 39
rect 25 36 29 39
rect -7 9 -3 32
rect 5 12 13 17
rect 25 9 29 32
rect -7 5 38 9
rect -21 -9 -6 -5
rect -21 -21 -17 -9
rect 1 -21 5 5
rect 13 -3 20 1
rect -55 -43 -45 -39
rect -55 -44 -51 -43
rect -63 -64 -59 -48
rect -29 -64 -25 -25
rect 9 -16 29 -12
rect 9 -21 13 -16
rect 25 -21 29 -16
rect -7 -32 -3 -27
rect 9 -32 13 -27
rect -7 -36 13 -32
rect -11 -43 4 -39
rect 17 -64 21 -27
rect -67 -68 -63 -64
rect -59 -68 37 -64
rect 41 -68 45 -64
<< metal2 >>
rect -66 12 -48 17
rect -71 3 -67 12
rect -38 1 -34 26
rect -25 12 1 17
rect -38 -3 9 1
rect -41 -43 -15 -39
<< ntransistor >>
rect -24 -25 -22 -21
rect -2 -28 0 -20
rect 6 -28 8 -20
rect 14 -28 16 -20
rect 22 -28 24 -20
rect -58 -48 -56 -44
<< ptransistor >>
rect -24 39 -22 49
rect -58 21 -56 31
rect -2 31 0 51
rect 6 31 8 51
rect 14 31 16 51
rect 22 31 24 51
<< polycontact >>
rect -28 26 -24 30
rect -62 -1 -58 3
rect -6 -9 -2 -5
rect 13 12 17 17
rect 20 -3 24 1
rect 4 -43 8 -39
<< ndcontact >>
rect -29 -25 -25 -21
rect -21 -25 -17 -21
rect -7 -27 -3 -21
rect 1 -27 5 -21
rect 9 -27 13 -21
rect 17 -27 21 -21
rect 25 -27 29 -21
rect -63 -48 -59 -44
rect -55 -48 -51 -44
<< pdcontact >>
rect -29 40 -25 48
rect -21 40 -17 48
rect -7 46 -3 50
rect -7 39 -3 43
rect -63 22 -59 30
rect -55 22 -51 30
rect -7 32 -3 36
rect 1 46 5 50
rect 1 39 5 43
rect 1 32 5 36
rect 9 46 13 50
rect 9 39 13 43
rect 9 32 13 36
rect 17 46 21 50
rect 17 39 21 43
rect 17 32 21 36
rect 25 46 29 50
rect 25 39 29 43
rect 25 32 29 36
<< m2contact >>
rect -38 26 -34 30
rect -71 12 -66 17
rect -71 -1 -67 3
rect -48 12 -43 17
rect -30 12 -25 17
rect 1 12 5 17
rect 9 -3 13 1
rect -45 -43 -41 -39
rect -15 -43 -11 -39
<< psubstratepcontact >>
rect -63 -68 -59 -64
rect 37 -68 41 -64
<< nsubstratencontact >>
rect -63 58 -59 62
rect 37 58 41 62
<< labels >>
rlabel nwell -67 58 45 62 0 Vdd
rlabel pwell -67 -68 45 -64 0 gnd
rlabel metal1 29 5 38 9 0 out
rlabel metal1 -75 -1 -71 3 0 b
rlabel metal1 -42 26 -38 30 0 a
<< end >>
