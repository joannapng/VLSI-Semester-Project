magic
tech scmos
timestamp 1672659533
<< polysilicon >>
rect -124 22 -22 24
rect -18 22 82 24
rect -124 14 -122 22
rect -32 6 -30 8
rect 80 6 82 22
rect -70 1 -68 3
rect -124 -4 -122 -2
rect 186 4 188 6
rect -124 -12 -122 -10
rect -124 -85 -122 -20
rect -93 -35 -91 -33
rect -93 -53 -91 -43
rect -70 -46 -68 -3
rect -56 -12 -54 -10
rect -32 -12 -30 -2
rect 80 -5 82 -2
rect 123 -6 145 -4
rect 80 -12 82 -9
rect -56 -21 -54 -16
rect -32 -18 -30 -16
rect -56 -45 -54 -25
rect -18 -26 -14 -24
rect 28 -28 30 -26
rect -18 -45 -14 -34
rect -70 -52 -68 -50
rect -18 -51 -14 -49
rect -93 -59 -91 -57
rect 28 -76 30 -32
rect 41 -37 43 -36
rect 41 -44 43 -41
rect 41 -56 43 -48
rect 28 -83 30 -80
rect 80 -85 82 -28
rect 123 -66 125 -6
rect 143 -9 145 -6
rect 143 -16 145 -13
rect 186 -14 188 -4
rect 186 -20 188 -18
rect 143 -23 145 -21
rect 200 -28 204 -26
rect 143 -35 145 -31
rect 143 -47 145 -39
rect 200 -47 204 -36
rect 248 -40 250 -38
rect 143 -54 145 -51
rect 200 -53 204 -51
rect 248 -58 250 -48
rect 143 -61 145 -59
rect 248 -64 250 -62
rect 123 -73 125 -70
rect 143 -73 145 -69
rect 123 -75 145 -73
rect -124 -87 -6 -85
rect -2 -87 82 -85
<< ndiffusion >>
rect -76 -3 -75 1
rect -71 -3 -70 1
rect -68 -3 -67 1
rect -63 -3 -62 1
rect 74 5 80 6
rect 74 -1 75 5
rect 79 -1 80 5
rect 74 -2 80 -1
rect 82 5 88 6
rect 82 -1 83 5
rect 87 -1 88 5
rect 82 -2 88 -1
rect -130 -13 -124 -12
rect -130 -19 -129 -13
rect -125 -19 -124 -13
rect -130 -20 -124 -19
rect -122 -13 -116 -12
rect -122 -19 -121 -13
rect -117 -19 -116 -13
rect -122 -20 -116 -19
rect -63 -16 -62 -12
rect -58 -16 -56 -12
rect -54 -16 -53 -12
rect -49 -16 -48 -12
rect -38 -16 -37 -12
rect -33 -16 -32 -12
rect -30 -16 -29 -12
rect -25 -16 -24 -12
rect 22 -32 23 -28
rect 27 -32 28 -28
rect 30 -32 31 -28
rect 35 -32 36 -28
rect -24 -49 -23 -45
rect -19 -49 -18 -45
rect -14 -49 -13 -45
rect -9 -49 -8 -45
rect -99 -57 -98 -53
rect -94 -57 -93 -53
rect -91 -57 -90 -53
rect -86 -57 -85 -53
rect 35 -48 36 -44
rect 40 -48 41 -44
rect 43 -48 44 -44
rect 48 -48 49 -44
rect 137 -13 138 -9
rect 142 -13 143 -9
rect 145 -13 146 -9
rect 150 -13 151 -9
rect 180 -18 181 -14
rect 185 -18 186 -14
rect 188 -18 189 -14
rect 193 -18 194 -14
rect 137 -51 138 -47
rect 142 -51 143 -47
rect 145 -51 146 -47
rect 150 -51 151 -47
rect 194 -51 195 -47
rect 199 -51 200 -47
rect 204 -51 205 -47
rect 209 -51 210 -47
rect 242 -62 243 -58
rect 247 -62 248 -58
rect 250 -62 251 -58
rect 255 -62 256 -58
<< pdiffusion >>
rect -130 13 -124 14
rect -130 -1 -129 13
rect -125 -1 -124 13
rect -130 -2 -124 -1
rect -122 13 -116 14
rect -122 -1 -121 13
rect -117 -1 -116 13
rect -38 5 -32 6
rect -122 -2 -116 -1
rect -38 -1 -37 5
rect -33 -1 -32 5
rect -38 -2 -32 -1
rect -30 5 -24 6
rect -30 -1 -29 5
rect -25 -1 -24 5
rect -30 -2 -24 -1
rect 180 3 186 4
rect -99 -36 -93 -35
rect -99 -42 -98 -36
rect -94 -42 -93 -36
rect -99 -43 -93 -42
rect -91 -36 -85 -35
rect -91 -42 -90 -36
rect -86 -42 -85 -36
rect -91 -43 -85 -42
rect 180 -3 181 3
rect 185 -3 186 3
rect 180 -4 186 -3
rect 188 3 194 4
rect 188 -3 189 3
rect 193 -3 194 3
rect 188 -4 194 -3
rect 74 -13 80 -12
rect -24 -27 -18 -26
rect -24 -33 -23 -27
rect -19 -33 -18 -27
rect -24 -34 -18 -33
rect -14 -27 -8 -26
rect -14 -33 -13 -27
rect -9 -33 -8 -27
rect 74 -27 75 -13
rect 79 -27 80 -13
rect 74 -28 80 -27
rect 82 -13 88 -12
rect 82 -27 83 -13
rect 87 -27 88 -13
rect 82 -28 88 -27
rect -14 -34 -8 -33
rect 137 -24 143 -23
rect 137 -30 138 -24
rect 142 -30 143 -24
rect 137 -31 143 -30
rect 145 -24 151 -23
rect 145 -30 146 -24
rect 150 -30 151 -24
rect 145 -31 151 -30
rect 194 -29 200 -28
rect 194 -35 195 -29
rect 199 -35 200 -29
rect 194 -36 200 -35
rect 204 -29 210 -28
rect 204 -35 205 -29
rect 209 -35 210 -29
rect 204 -36 210 -35
rect 242 -41 248 -40
rect 242 -47 243 -41
rect 247 -47 248 -41
rect 242 -48 248 -47
rect 250 -41 256 -40
rect 250 -47 251 -41
rect 255 -47 256 -41
rect 250 -48 256 -47
rect 137 -62 143 -61
rect 137 -68 138 -62
rect 142 -68 143 -62
rect 137 -69 143 -68
rect 145 -62 151 -61
rect 145 -68 146 -62
rect 150 -68 151 -62
rect 145 -69 151 -68
<< metal1 >>
rect -131 31 247 35
rect -98 17 -94 31
rect -129 -5 -125 -1
rect -135 -9 -125 -5
rect -129 -13 -125 -9
rect -37 5 -33 31
rect -13 7 -9 31
rect -121 -5 -117 -1
rect -110 -3 -75 1
rect -63 -3 -49 1
rect 63 9 114 13
rect -110 -5 -106 -3
rect -121 -9 -106 -5
rect -53 -5 -49 -3
rect -29 -5 -25 -1
rect 63 -5 68 9
rect 75 -5 79 -1
rect -53 -9 -36 -5
rect -29 -9 79 -5
rect -121 -13 -117 -9
rect -114 -30 -110 -9
rect -53 -12 -49 -9
rect -29 -12 -25 -9
rect -78 -16 -62 -12
rect -78 -21 -74 -16
rect -105 -25 -57 -21
rect -105 -46 -101 -25
rect -98 -36 -94 -32
rect -90 -46 -86 -42
rect -107 -50 -97 -46
rect -90 -50 -71 -46
rect -90 -53 -86 -50
rect -98 -92 -94 -57
rect -80 -76 -76 -50
rect -64 -66 -60 -25
rect -37 -92 -33 -16
rect -13 -27 -9 -23
rect 46 -28 50 -9
rect 75 -13 79 -9
rect 83 -5 87 -1
rect 83 -9 99 -5
rect 83 -13 87 -9
rect 95 -24 99 -9
rect 110 -16 114 9
rect 181 3 185 31
rect 205 5 209 31
rect 189 -7 193 -3
rect 138 -16 142 -13
rect 110 -20 142 -16
rect 138 -24 142 -20
rect 16 -32 23 -28
rect 35 -32 50 -28
rect 95 -28 107 -24
rect -23 -37 -19 -33
rect 16 -37 20 -32
rect -24 -41 -19 -37
rect -10 -41 20 -37
rect 37 -41 41 -37
rect -23 -45 -19 -41
rect 16 -44 20 -41
rect 16 -48 36 -44
rect 40 -48 41 -44
rect -13 -92 -9 -49
rect 44 -59 48 -48
rect 95 -54 99 -28
rect 146 -16 150 -13
rect 162 -11 182 -7
rect 189 -11 234 -7
rect 162 -16 166 -11
rect 189 -14 193 -11
rect 146 -20 166 -16
rect 146 -24 150 -20
rect 110 -39 142 -35
rect 138 -54 142 -51
rect 15 -63 48 -59
rect 95 -58 142 -54
rect 15 -69 19 -63
rect 56 -69 60 -59
rect 138 -62 142 -58
rect 15 -73 60 -69
rect 109 -70 122 -66
rect 146 -54 150 -51
rect 155 -54 159 -20
rect 146 -58 159 -54
rect 146 -62 150 -58
rect 15 -76 19 -73
rect 11 -80 27 -76
rect 181 -92 185 -18
rect 205 -29 209 -25
rect 195 -39 199 -35
rect 214 -39 218 -11
rect 194 -43 199 -39
rect 208 -43 218 -39
rect 195 -47 199 -43
rect 205 -92 209 -51
rect 230 -51 234 -11
rect 243 -41 247 31
rect 251 -51 255 -47
rect 230 -55 244 -51
rect 251 -55 263 -51
rect 251 -58 255 -55
rect 243 -92 247 -62
rect -127 -96 247 -92
<< metal2 >>
rect -98 -28 -94 13
rect -13 -19 -9 3
rect 205 -21 209 1
rect 111 -28 123 -24
rect -114 -37 -110 -34
rect -114 -41 -28 -37
rect -4 -41 33 -37
rect -4 -66 0 -41
rect 106 -55 110 -39
rect 119 -39 123 -28
rect 119 -43 190 -39
rect 60 -59 110 -55
rect -60 -70 105 -66
rect -76 -80 7 -76
<< ntransistor >>
rect -70 -3 -68 1
rect 80 -2 82 6
rect -124 -20 -122 -12
rect -56 -16 -54 -12
rect -32 -16 -30 -12
rect 28 -32 30 -28
rect -18 -49 -14 -45
rect -93 -57 -91 -53
rect 41 -48 43 -44
rect 143 -13 145 -9
rect 186 -18 188 -14
rect 143 -51 145 -47
rect 200 -51 204 -47
rect 248 -62 250 -58
<< ptransistor >>
rect -124 -2 -122 14
rect -32 -2 -30 6
rect -93 -43 -91 -35
rect 186 -4 188 4
rect -18 -34 -14 -26
rect 80 -28 82 -12
rect 143 -31 145 -23
rect 200 -36 204 -28
rect 248 -48 250 -40
rect 143 -69 145 -61
<< polycontact >>
rect -22 22 -18 26
rect -97 -50 -93 -46
rect -36 -9 -32 -5
rect -57 -25 -53 -21
rect -14 -41 -10 -37
rect -71 -50 -67 -46
rect 41 -41 45 -37
rect 27 -80 31 -76
rect 182 -11 186 -7
rect 142 -39 146 -35
rect 204 -43 208 -39
rect 244 -55 248 -51
rect 122 -70 126 -66
rect -6 -89 -2 -85
<< ndcontact >>
rect -75 -3 -71 1
rect -67 -3 -63 1
rect 75 -1 79 5
rect 83 -1 87 5
rect -129 -19 -125 -13
rect -121 -19 -117 -13
rect -62 -16 -58 -12
rect -53 -16 -49 -12
rect -37 -16 -33 -12
rect -29 -16 -25 -12
rect 23 -32 27 -28
rect 31 -32 35 -28
rect -23 -49 -19 -45
rect -13 -49 -9 -45
rect -98 -57 -94 -53
rect -90 -57 -86 -53
rect 36 -48 40 -44
rect 44 -48 48 -44
rect 138 -13 142 -9
rect 146 -13 150 -9
rect 181 -18 185 -14
rect 189 -18 193 -14
rect 138 -51 142 -47
rect 146 -51 150 -47
rect 195 -51 199 -47
rect 205 -51 209 -47
rect 243 -62 247 -58
rect 251 -62 255 -58
<< pdcontact >>
rect -129 -1 -125 13
rect -121 -1 -117 13
rect -37 -1 -33 5
rect -29 -1 -25 5
rect -98 -42 -94 -36
rect -90 -42 -86 -36
rect 181 -3 185 3
rect 189 -3 193 3
rect -23 -33 -19 -27
rect -13 -33 -9 -27
rect 75 -27 79 -13
rect 83 -27 87 -13
rect 138 -30 142 -24
rect 146 -30 150 -24
rect 195 -35 199 -29
rect 205 -35 209 -29
rect 243 -47 247 -41
rect 251 -47 255 -41
rect 138 -68 142 -62
rect 146 -68 150 -62
<< m2contact >>
rect -98 13 -94 17
rect -13 3 -9 7
rect -114 -34 -110 -30
rect -98 -32 -94 -28
rect -64 -70 -60 -66
rect -80 -80 -76 -76
rect -13 -23 -9 -19
rect 205 1 209 5
rect 107 -28 111 -24
rect -28 -41 -24 -37
rect 33 -41 37 -37
rect 106 -39 110 -35
rect 56 -59 60 -55
rect 105 -70 109 -66
rect 7 -80 11 -76
rect 205 -25 209 -21
rect 190 -43 194 -39
<< labels >>
rlabel metal1 -135 -9 -129 -5 0 D
rlabel polycontact -22 22 -18 26 0 clk
rlabel metal1 -107 -50 -99 -46 0 S
rlabel metal1 49 -9 56 -5 0 Qm
rlabel metal1 -131 31 209 35 0 Vdd
rlabel metal1 87 -9 99 -5 0 Qpass
rlabel metal1 154 -20 166 -16 1 mux_out_1
rlabel polycontact -6 -89 -2 -85 0 not_clk
rlabel metal1 -114 -9 -106 -5 0 Dpass
rlabel metal1 218 -11 230 -7 0 Q
rlabel metal1 -49 -9 -40 -5 0 or_1_out
rlabel metal1 -10 -41 -4 -37 0 or_2_out
rlabel metal1 -90 -50 -79 -46 0 not_S
rlabel metal1 -127 -96 209 -92 0 gnd
rlabel metal1 255 -55 263 -51 0 Qbar
<< end >>
