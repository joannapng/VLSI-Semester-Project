.include "d_ff_async_set_reset.spice"

.param vdd=2.5V clk_period=20u half_period=10u tr=10p tf=10p td=10u wnmin=3u wpmin=9u


Vdd Vdd 0 DC vdd
Vclk clk 0 pulse (0 {vdd} {td} {tr} {tf} {half_period} {clk_period})
Vnot_clk not_clk 0 pulse (0 {vdd} 0 {tr} {tf} {half_period} {clk_period})

Vs S 0 pwl (
    + 0 0 
    + 3u 0
    + {3u + 10p} {vdd}
    + 8u {vdd}
    + {8u + 10p} 0
    + 45u   0
    + {45u+10p} {vdd}
    + 55u   {vdd}
    + {55u + 10p} 0
+)

Vr R 0 pwl (
    + 0 0 
    + 23u 0
    + {23u + 10p} {vdd}
    + 28u {vdd}
    + {28u + 10p} 0
    + 53u 0
    + {53u+10p} {vdd}
    + 65u {vdd}
    + {65u+10p} 0
+)

Vd D 0 pwl (
    + 0 0 
    + 6u 0
    + {6u + 10p} {vdd}
    + 24u {vdd}
    + {24u + 10p} 0
    + 28u   0
    + {28u+10p} {vdd}
    + 34u {vdd}
    + {34u+10p} {0}
    + 68u   {0}
    + {68u +10p} {vdd}
    + 75u       {vdd}
    + {75u + 10p} 0
+)

.ic V(Q)=0
.tran 100n 110u

.control
    run
    set xbrushwidth=3
    set color0=white
    set color1=black
    set hcopyheight=200
    set hcopywidth=1000
    set hcopydevtype=svg
.endc

.end
