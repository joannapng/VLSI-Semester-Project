magic
tech scmos
timestamp 1672503769
<< polysilicon >>
rect -6 22 27 24
rect 31 22 63 24
rect -6 6 -4 22
rect 17 6 19 8
rect 61 2 63 22
rect 86 6 88 8
rect -6 -4 -4 -2
rect -6 -12 -4 -10
rect 17 -12 19 -2
rect 61 -5 63 -2
rect 61 -12 63 -9
rect 86 -12 88 -2
rect 137 -12 139 -10
rect -6 -63 -4 -16
rect 17 -18 19 -16
rect 86 -18 88 -16
rect 31 -26 35 -24
rect 31 -45 35 -34
rect 31 -51 35 -49
rect 61 -63 63 -20
rect 100 -26 104 -24
rect 137 -30 139 -20
rect 100 -45 104 -34
rect 137 -36 139 -34
rect 100 -51 104 -49
rect -6 -65 43 -63
rect 47 -65 63 -63
<< ndiffusion >>
rect 55 -2 56 2
rect 60 -2 61 2
rect 63 -2 64 2
rect 68 -2 69 2
rect -12 -16 -11 -12
rect -7 -16 -6 -12
rect -4 -16 -3 -12
rect 1 -16 2 -12
rect 11 -16 12 -12
rect 16 -16 17 -12
rect 19 -16 20 -12
rect 24 -16 25 -12
rect 80 -16 81 -12
rect 85 -16 86 -12
rect 88 -16 89 -12
rect 93 -16 94 -12
rect 25 -49 26 -45
rect 30 -49 31 -45
rect 35 -49 36 -45
rect 40 -49 41 -45
rect 131 -34 132 -30
rect 136 -34 137 -30
rect 139 -34 140 -30
rect 144 -34 145 -30
rect 94 -49 95 -45
rect 99 -49 100 -45
rect 104 -49 105 -45
rect 109 -49 110 -45
<< pdiffusion >>
rect -12 5 -6 6
rect -12 -1 -11 5
rect -7 -1 -6 5
rect -12 -2 -6 -1
rect -4 5 2 6
rect -4 -1 -3 5
rect 1 -1 2 5
rect -4 -2 2 -1
rect 11 5 17 6
rect 11 -1 12 5
rect 16 -1 17 5
rect 11 -2 17 -1
rect 19 5 25 6
rect 19 -1 20 5
rect 24 -1 25 5
rect 80 5 86 6
rect 19 -2 25 -1
rect 80 -1 81 5
rect 85 -1 86 5
rect 80 -2 86 -1
rect 88 5 94 6
rect 88 -1 89 5
rect 93 -1 94 5
rect 88 -2 94 -1
rect 55 -13 61 -12
rect 55 -19 56 -13
rect 60 -19 61 -13
rect 55 -20 61 -19
rect 63 -13 69 -12
rect 63 -19 64 -13
rect 68 -19 69 -13
rect 131 -13 137 -12
rect 63 -20 69 -19
rect 131 -19 132 -13
rect 136 -19 137 -13
rect 131 -20 137 -19
rect 139 -13 145 -12
rect 139 -19 140 -13
rect 144 -19 145 -13
rect 139 -20 145 -19
rect 25 -27 31 -26
rect 25 -33 26 -27
rect 30 -33 31 -27
rect 25 -34 31 -33
rect 35 -27 41 -26
rect 35 -33 36 -27
rect 40 -33 41 -27
rect 35 -34 41 -33
rect 94 -27 100 -26
rect 94 -33 95 -27
rect 99 -33 100 -27
rect 94 -34 100 -33
rect 104 -27 110 -26
rect 104 -33 105 -27
rect 109 -33 110 -27
rect 104 -34 110 -33
<< metal1 >>
rect -13 31 136 35
rect 12 5 16 31
rect 36 7 40 31
rect -11 -5 -7 -1
rect -17 -9 -7 -5
rect -11 -12 -7 -9
rect 81 5 85 31
rect 105 7 109 31
rect -3 -5 1 -1
rect 20 -5 24 -1
rect 56 -5 60 -2
rect -3 -9 13 -5
rect 20 -9 60 -5
rect -3 -12 1 -9
rect 4 -30 8 -9
rect 20 -12 24 -9
rect 12 -70 16 -16
rect 36 -27 40 -23
rect 26 -37 30 -33
rect 45 -37 49 -9
rect 56 -13 60 -9
rect 64 -5 68 -2
rect 89 -5 93 -1
rect 64 -9 82 -5
rect 89 -9 128 -5
rect 64 -13 68 -9
rect 73 -30 77 -9
rect 89 -12 93 -9
rect 25 -41 30 -37
rect 39 -41 49 -37
rect 26 -45 30 -41
rect 36 -70 40 -49
rect 81 -70 85 -16
rect 105 -27 109 -23
rect 95 -37 99 -33
rect 114 -37 118 -9
rect 124 -23 128 -9
rect 132 -13 136 31
rect 140 -23 144 -19
rect 124 -27 133 -23
rect 140 -27 153 -23
rect 140 -30 144 -27
rect 94 -41 99 -37
rect 108 -41 118 -37
rect 95 -45 99 -41
rect 105 -70 109 -49
rect 132 -70 136 -34
rect -13 -74 136 -70
<< metal2 >>
rect 36 -19 40 3
rect 105 -19 109 3
rect 4 -37 8 -34
rect 73 -37 77 -34
rect 4 -41 21 -37
rect 73 -41 90 -37
<< ntransistor >>
rect 61 -2 63 2
rect -6 -16 -4 -12
rect 17 -16 19 -12
rect 86 -16 88 -12
rect 31 -49 35 -45
rect 137 -34 139 -30
rect 100 -49 104 -45
<< ptransistor >>
rect -6 -2 -4 6
rect 17 -2 19 6
rect 86 -2 88 6
rect 61 -20 63 -12
rect 137 -20 139 -12
rect 31 -34 35 -26
rect 100 -34 104 -26
<< polycontact >>
rect 27 22 31 26
rect 13 -9 17 -5
rect 82 -9 86 -5
rect 35 -41 39 -37
rect 133 -27 137 -23
rect 104 -41 108 -37
rect 43 -67 47 -63
<< ndcontact >>
rect 56 -2 60 2
rect 64 -2 68 2
rect -11 -16 -7 -12
rect -3 -16 1 -12
rect 12 -16 16 -12
rect 20 -16 24 -12
rect 81 -16 85 -12
rect 89 -16 93 -12
rect 26 -49 30 -45
rect 36 -49 40 -45
rect 132 -34 136 -30
rect 140 -34 144 -30
rect 95 -49 99 -45
rect 105 -49 109 -45
<< pdcontact >>
rect -11 -1 -7 5
rect -3 -1 1 5
rect 12 -1 16 5
rect 20 -1 24 5
rect 81 -1 85 5
rect 89 -1 93 5
rect 56 -19 60 -13
rect 64 -19 68 -13
rect 132 -19 136 -13
rect 140 -19 144 -13
rect 26 -33 30 -27
rect 36 -33 40 -27
rect 95 -33 99 -27
rect 105 -33 109 -27
<< m2contact >>
rect 36 3 40 7
rect 4 -34 8 -30
rect 36 -23 40 -19
rect 105 3 109 7
rect 73 -34 77 -30
rect 21 -41 25 -37
rect 105 -23 109 -19
rect 90 -41 94 -37
<< labels >>
rlabel polycontact 27 22 31 26 0 clk
rlabel metal1 49 -9 56 -5 0 Qm
rlabel metal1 112 -9 121 -5 0 Q
rlabel polycontact 43 -67 47 -63 0 not_clk
rlabel metal1 -17 -9 -11 -5 0 D
rlabel metal1 144 -27 153 -23 0 Qbar
rlabel metal1 -13 31 136 35 0 Vdd
rlabel metal1 -13 -74 136 -70 0 gnd
<< end >>
