magic
tech scmos
timestamp 1671962531
<< polysilicon >>
rect -124 22 -22 24
rect -18 22 63 24
rect -124 14 -122 22
rect -32 6 -30 8
rect 61 6 63 22
rect 86 6 88 8
rect -70 1 -68 3
rect -124 -4 -122 -2
rect -124 -12 -122 -10
rect -124 -85 -122 -20
rect -93 -35 -91 -33
rect -93 -53 -91 -43
rect -70 -46 -68 -3
rect -56 -12 -54 -10
rect -32 -12 -30 -2
rect 61 -5 63 -2
rect 61 -12 63 -9
rect 86 -12 88 -2
rect -56 -21 -54 -16
rect -32 -18 -30 -16
rect -56 -45 -54 -25
rect -18 -26 -14 -24
rect 28 -28 30 -26
rect 86 -18 88 -16
rect 100 -26 104 -24
rect -18 -45 -14 -34
rect -70 -52 -68 -50
rect -18 -51 -14 -49
rect -93 -59 -91 -57
rect 28 -76 30 -32
rect 41 -37 43 -36
rect 41 -44 43 -41
rect 41 -56 43 -48
rect 28 -85 30 -80
rect 61 -85 63 -28
rect 100 -45 104 -34
rect 100 -51 104 -49
rect -124 -87 -6 -85
rect -2 -87 63 -85
<< ndiffusion >>
rect -76 -3 -75 1
rect -71 -3 -70 1
rect -68 -3 -67 1
rect -63 -3 -62 1
rect 55 5 61 6
rect 55 -1 56 5
rect 60 -1 61 5
rect 55 -2 61 -1
rect 63 5 69 6
rect 63 -1 64 5
rect 68 -1 69 5
rect 63 -2 69 -1
rect -130 -13 -124 -12
rect -130 -19 -129 -13
rect -125 -19 -124 -13
rect -130 -20 -124 -19
rect -122 -13 -116 -12
rect -122 -19 -121 -13
rect -117 -19 -116 -13
rect -122 -20 -116 -19
rect -63 -16 -62 -12
rect -58 -16 -56 -12
rect -54 -16 -53 -12
rect -49 -16 -48 -12
rect -38 -16 -37 -12
rect -33 -16 -32 -12
rect -30 -16 -29 -12
rect -25 -16 -24 -12
rect 80 -16 81 -12
rect 85 -16 86 -12
rect 88 -16 89 -12
rect 93 -16 94 -12
rect 22 -32 23 -28
rect 27 -32 28 -28
rect 30 -32 31 -28
rect 35 -32 36 -28
rect -24 -49 -23 -45
rect -19 -49 -18 -45
rect -14 -49 -13 -45
rect -9 -49 -8 -45
rect -99 -57 -98 -53
rect -94 -57 -93 -53
rect -91 -57 -90 -53
rect -86 -57 -85 -53
rect 35 -48 36 -44
rect 40 -48 41 -44
rect 43 -48 44 -44
rect 48 -48 49 -44
rect 94 -49 95 -45
rect 99 -49 100 -45
rect 104 -49 105 -45
rect 109 -49 110 -45
<< pdiffusion >>
rect -130 13 -124 14
rect -130 -1 -129 13
rect -125 -1 -124 13
rect -130 -2 -124 -1
rect -122 13 -116 14
rect -122 -1 -121 13
rect -117 -1 -116 13
rect -38 5 -32 6
rect -122 -2 -116 -1
rect -38 -1 -37 5
rect -33 -1 -32 5
rect -38 -2 -32 -1
rect -30 5 -24 6
rect -30 -1 -29 5
rect -25 -1 -24 5
rect -30 -2 -24 -1
rect 80 5 86 6
rect 80 -1 81 5
rect 85 -1 86 5
rect 80 -2 86 -1
rect 88 5 94 6
rect 88 -1 89 5
rect 93 -1 94 5
rect 88 -2 94 -1
rect -99 -36 -93 -35
rect -99 -42 -98 -36
rect -94 -42 -93 -36
rect -99 -43 -93 -42
rect -91 -36 -85 -35
rect -91 -42 -90 -36
rect -86 -42 -85 -36
rect -91 -43 -85 -42
rect 55 -13 61 -12
rect -24 -27 -18 -26
rect -24 -33 -23 -27
rect -19 -33 -18 -27
rect -24 -34 -18 -33
rect -14 -27 -8 -26
rect -14 -33 -13 -27
rect -9 -33 -8 -27
rect 55 -27 56 -13
rect 60 -27 61 -13
rect 55 -28 61 -27
rect 63 -13 69 -12
rect 63 -27 64 -13
rect 68 -27 69 -13
rect 63 -28 69 -27
rect 94 -27 100 -26
rect -14 -34 -8 -33
rect 94 -33 95 -27
rect 99 -33 100 -27
rect 94 -34 100 -33
rect 104 -27 110 -26
rect 104 -33 105 -27
rect 109 -33 110 -27
rect 104 -34 110 -33
<< metal1 >>
rect -131 31 109 35
rect -98 17 -94 31
rect -129 -5 -125 -1
rect -135 -9 -125 -5
rect -129 -13 -125 -9
rect -37 5 -33 31
rect -13 7 -9 31
rect -121 -5 -117 -1
rect -110 -3 -75 1
rect -63 -3 -49 1
rect 81 5 85 31
rect 105 7 109 31
rect -110 -5 -106 -3
rect -121 -9 -106 -5
rect -53 -5 -49 -3
rect -29 -5 -25 -1
rect 56 -5 60 -1
rect -53 -9 -36 -5
rect -29 -9 60 -5
rect -121 -13 -117 -9
rect -114 -30 -110 -9
rect -53 -12 -49 -9
rect -29 -12 -25 -9
rect -78 -16 -62 -12
rect -78 -21 -74 -16
rect -105 -25 -57 -21
rect -105 -46 -101 -25
rect -98 -36 -94 -32
rect -90 -46 -86 -42
rect -107 -50 -97 -46
rect -90 -50 -71 -46
rect -90 -53 -86 -50
rect -98 -92 -94 -57
rect -80 -76 -76 -50
rect -64 -66 -60 -25
rect -37 -92 -33 -16
rect -13 -27 -9 -23
rect 46 -28 50 -9
rect 56 -13 60 -9
rect 64 -5 68 -1
rect 89 -5 93 -1
rect 64 -9 82 -5
rect 89 -9 121 -5
rect 64 -13 68 -9
rect 16 -32 23 -28
rect 35 -32 50 -28
rect 73 -30 77 -9
rect 89 -12 93 -9
rect -23 -37 -19 -33
rect 16 -37 20 -32
rect -24 -41 -19 -37
rect -10 -41 20 -37
rect 37 -41 41 -37
rect -23 -45 -19 -41
rect 16 -44 20 -41
rect 16 -48 36 -44
rect 40 -48 41 -44
rect -13 -92 -9 -49
rect 44 -63 48 -48
rect 15 -67 48 -63
rect 15 -76 19 -67
rect 11 -80 27 -76
rect 81 -92 85 -16
rect 105 -27 109 -23
rect 95 -37 99 -33
rect 114 -37 118 -9
rect 94 -41 99 -37
rect 108 -41 118 -37
rect 95 -45 99 -41
rect 105 -92 109 -49
rect -131 -96 109 -92
<< metal2 >>
rect -98 -28 -94 13
rect -13 -19 -9 3
rect 105 -19 109 3
rect -114 -37 -110 -34
rect 73 -37 77 -34
rect -114 -41 -28 -37
rect -4 -41 33 -37
rect 73 -41 90 -37
rect -4 -66 0 -41
rect -60 -70 0 -66
rect -76 -80 7 -76
<< ntransistor >>
rect -70 -3 -68 1
rect 61 -2 63 6
rect -124 -20 -122 -12
rect -56 -16 -54 -12
rect -32 -16 -30 -12
rect 86 -16 88 -12
rect 28 -32 30 -28
rect -18 -49 -14 -45
rect -93 -57 -91 -53
rect 41 -48 43 -44
rect 100 -49 104 -45
<< ptransistor >>
rect -124 -2 -122 14
rect -32 -2 -30 6
rect 86 -2 88 6
rect -93 -43 -91 -35
rect -18 -34 -14 -26
rect 61 -28 63 -12
rect 100 -34 104 -26
<< polycontact >>
rect -22 22 -18 26
rect -97 -50 -93 -46
rect -36 -9 -32 -5
rect 82 -9 86 -5
rect -57 -25 -53 -21
rect -14 -41 -10 -37
rect -71 -50 -67 -46
rect 41 -41 45 -37
rect 27 -80 31 -76
rect 104 -41 108 -37
rect -6 -89 -2 -85
<< ndcontact >>
rect -75 -3 -71 1
rect -67 -3 -63 1
rect 56 -1 60 5
rect 64 -1 68 5
rect -129 -19 -125 -13
rect -121 -19 -117 -13
rect -62 -16 -58 -12
rect -53 -16 -49 -12
rect -37 -16 -33 -12
rect -29 -16 -25 -12
rect 81 -16 85 -12
rect 89 -16 93 -12
rect 23 -32 27 -28
rect 31 -32 35 -28
rect -23 -49 -19 -45
rect -13 -49 -9 -45
rect -98 -57 -94 -53
rect -90 -57 -86 -53
rect 36 -48 40 -44
rect 44 -48 48 -44
rect 95 -49 99 -45
rect 105 -49 109 -45
<< pdcontact >>
rect -129 -1 -125 13
rect -121 -1 -117 13
rect -37 -1 -33 5
rect -29 -1 -25 5
rect 81 -1 85 5
rect 89 -1 93 5
rect -98 -42 -94 -36
rect -90 -42 -86 -36
rect -23 -33 -19 -27
rect -13 -33 -9 -27
rect 56 -27 60 -13
rect 64 -27 68 -13
rect 95 -33 99 -27
rect 105 -33 109 -27
<< m2contact >>
rect -98 13 -94 17
rect -13 3 -9 7
rect -114 -34 -110 -30
rect -98 -32 -94 -28
rect -64 -70 -60 -66
rect -80 -80 -76 -76
rect -13 -23 -9 -19
rect 105 3 109 7
rect 73 -34 77 -30
rect -28 -41 -24 -37
rect 33 -41 37 -37
rect 7 -80 11 -76
rect 105 -23 109 -19
rect 90 -41 94 -37
<< labels >>
rlabel metal1 49 -9 56 -5 0 Qm
rlabel metal1 112 -9 121 -5 0 Q
rlabel metal1 -135 -9 -129 -5 0 D
rlabel polycontact -22 22 -18 26 0 clk
rlabel metal1 -107 -50 -99 -46 0 S
rlabel polycontact -6 -89 -2 -85 0 not_clk
rlabel metal1 -131 31 109 35 0 Vdd
rlabel metal1 -131 -96 109 -92 0 gnd
<< end >>
