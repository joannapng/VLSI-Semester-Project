magic
tech scmos
timestamp 1671461162
<< polysilicon >>
rect 267 39 269 44
rect 267 32 269 35
rect 267 30 293 32
rect 152 28 154 30
rect 172 28 200 30
rect 267 28 269 30
rect -6 22 27 24
rect 31 22 63 24
rect -6 14 -4 22
rect 17 6 19 8
rect 61 6 63 22
rect 152 10 154 20
rect 172 17 174 28
rect 198 22 200 28
rect 267 18 269 20
rect 86 6 88 8
rect 152 4 154 6
rect -6 -4 -4 -2
rect -6 -12 -4 -10
rect 17 -12 19 -2
rect 61 -5 63 -2
rect 61 -12 63 -9
rect 86 -12 88 -2
rect 17 -18 19 -16
rect -6 -63 -4 -20
rect 31 -26 35 -24
rect 86 -18 88 -16
rect 100 -26 104 -24
rect 31 -45 35 -34
rect 31 -51 35 -49
rect 61 -63 63 -28
rect 100 -45 104 -34
rect 172 -43 174 13
rect 198 12 200 14
rect 267 9 269 11
rect 198 3 200 5
rect 198 -5 200 -3
rect 245 -8 247 -6
rect 198 -15 200 -9
rect 198 -25 200 -23
rect 245 -26 247 -16
rect 267 -19 269 3
rect 245 -32 247 -30
rect 198 -34 200 -32
rect 198 -43 200 -40
rect 267 -42 269 -23
rect 172 -45 200 -43
rect 100 -51 104 -49
rect 267 -52 269 -50
rect 267 -61 269 -59
rect -6 -65 43 -63
rect 47 -65 63 -63
rect 267 -69 269 -67
rect 291 -69 293 30
rect 267 -71 293 -69
<< ndiffusion >>
rect 146 6 147 10
rect 151 6 152 10
rect 154 6 155 10
rect 159 6 160 10
rect 55 5 61 6
rect 55 -1 56 5
rect 60 -1 61 5
rect 55 -2 61 -1
rect 63 5 69 6
rect 63 -1 64 5
rect 68 -1 69 5
rect 63 -2 69 -1
rect -12 -13 -6 -12
rect -12 -19 -11 -13
rect -7 -19 -6 -13
rect -12 -20 -6 -19
rect -4 -13 2 -12
rect -4 -19 -3 -13
rect 1 -19 2 -13
rect 11 -16 12 -12
rect 16 -16 17 -12
rect 19 -16 20 -12
rect 24 -16 25 -12
rect -4 -20 2 -19
rect 80 -16 81 -12
rect 85 -16 86 -12
rect 88 -16 89 -12
rect 93 -16 94 -12
rect 25 -49 26 -45
rect 30 -49 31 -45
rect 35 -49 36 -45
rect 40 -49 41 -45
rect 261 8 267 9
rect 261 4 262 8
rect 266 4 267 8
rect 261 3 267 4
rect 269 8 275 9
rect 269 4 270 8
rect 274 4 275 8
rect 269 3 275 4
rect 192 2 198 3
rect 192 -2 193 2
rect 197 -2 198 2
rect 192 -3 198 -2
rect 200 2 206 3
rect 200 -2 201 2
rect 205 -2 206 2
rect 200 -3 206 -2
rect 239 -30 240 -26
rect 244 -30 245 -26
rect 247 -30 248 -26
rect 252 -30 253 -26
rect 192 -35 198 -34
rect 192 -39 193 -35
rect 197 -39 198 -35
rect 192 -40 198 -39
rect 200 -35 206 -34
rect 200 -39 201 -35
rect 205 -39 206 -35
rect 200 -40 206 -39
rect 94 -49 95 -45
rect 99 -49 100 -45
rect 104 -49 105 -45
rect 109 -49 110 -45
rect 261 -62 267 -61
rect 261 -66 262 -62
rect 266 -66 267 -62
rect 261 -67 267 -66
rect 269 -62 275 -61
rect 269 -66 270 -62
rect 274 -66 275 -62
rect 269 -67 275 -66
<< pdiffusion >>
rect 146 27 152 28
rect -12 13 -6 14
rect -12 -1 -11 13
rect -7 -1 -6 13
rect -12 -2 -6 -1
rect -4 13 2 14
rect -4 -1 -3 13
rect 1 -1 2 13
rect 146 21 147 27
rect 151 21 152 27
rect 146 20 152 21
rect 154 27 160 28
rect 154 21 155 27
rect 159 21 160 27
rect 154 20 160 21
rect 261 27 267 28
rect 192 21 198 22
rect 192 15 193 21
rect 197 15 198 21
rect 192 14 198 15
rect 200 21 206 22
rect 200 15 201 21
rect 205 15 206 21
rect 261 21 262 27
rect 266 21 267 27
rect 261 20 267 21
rect 269 27 275 28
rect 269 21 270 27
rect 274 21 275 27
rect 269 20 275 21
rect 200 14 206 15
rect -4 -2 2 -1
rect 11 5 17 6
rect 11 -1 12 5
rect 16 -1 17 5
rect 11 -2 17 -1
rect 19 5 25 6
rect 19 -1 20 5
rect 24 -1 25 5
rect 19 -2 25 -1
rect 80 5 86 6
rect 80 -1 81 5
rect 85 -1 86 5
rect 80 -2 86 -1
rect 88 5 94 6
rect 88 -1 89 5
rect 93 -1 94 5
rect 88 -2 94 -1
rect 55 -13 61 -12
rect 25 -27 31 -26
rect 25 -33 26 -27
rect 30 -33 31 -27
rect 25 -34 31 -33
rect 35 -27 41 -26
rect 35 -33 36 -27
rect 40 -33 41 -27
rect 55 -27 56 -13
rect 60 -27 61 -13
rect 55 -28 61 -27
rect 63 -13 69 -12
rect 63 -27 64 -13
rect 68 -27 69 -13
rect 63 -28 69 -27
rect 94 -27 100 -26
rect 35 -34 41 -33
rect 94 -33 95 -27
rect 99 -33 100 -27
rect 94 -34 100 -33
rect 104 -27 110 -26
rect 104 -33 105 -27
rect 109 -33 110 -27
rect 104 -34 110 -33
rect 239 -9 245 -8
rect 239 -15 240 -9
rect 244 -15 245 -9
rect 192 -16 198 -15
rect 192 -22 193 -16
rect 197 -22 198 -16
rect 192 -23 198 -22
rect 200 -16 206 -15
rect 239 -16 245 -15
rect 247 -9 253 -8
rect 247 -15 248 -9
rect 252 -15 253 -9
rect 247 -16 253 -15
rect 200 -22 201 -16
rect 205 -22 206 -16
rect 200 -23 206 -22
rect 261 -43 267 -42
rect 261 -49 262 -43
rect 266 -49 267 -43
rect 261 -50 267 -49
rect 269 -43 275 -42
rect 269 -49 270 -43
rect 274 -49 275 -43
rect 269 -50 275 -49
<< metal1 >>
rect 229 35 265 39
rect -16 31 189 35
rect -11 -5 -7 -1
rect -25 -10 -7 -5
rect -11 -13 -7 -10
rect 12 5 16 31
rect 36 7 40 31
rect 81 5 85 31
rect 105 7 109 31
rect 147 27 151 31
rect 155 17 159 21
rect -3 -5 1 -1
rect 20 -5 24 -1
rect 56 -5 60 -1
rect -3 -9 13 -5
rect 20 -9 60 -5
rect -3 -13 1 -9
rect 4 -30 8 -9
rect 20 -12 24 -9
rect 12 -70 16 -16
rect 36 -27 40 -23
rect 26 -37 30 -33
rect 45 -37 49 -9
rect 56 -13 60 -9
rect 132 13 148 17
rect 155 13 170 17
rect 64 -5 68 -1
rect 89 -5 93 -1
rect 132 -5 136 13
rect 155 10 159 13
rect 185 10 189 31
rect 193 10 197 15
rect 185 6 197 10
rect 147 4 151 6
rect 193 2 197 6
rect 262 16 266 21
rect 201 11 205 15
rect 252 12 266 16
rect 201 7 213 11
rect 201 2 205 7
rect 209 -1 213 7
rect 252 -1 256 12
rect 262 8 266 12
rect 270 17 274 21
rect 270 13 282 17
rect 270 8 274 13
rect 209 -5 256 -1
rect 64 -9 82 -5
rect 89 -9 127 -5
rect 132 -9 196 -5
rect 64 -13 68 -9
rect 73 -30 77 -9
rect 89 -12 93 -9
rect 25 -41 30 -37
rect 39 -41 49 -37
rect 26 -45 30 -41
rect 36 -70 40 -49
rect 81 -70 85 -16
rect 105 -27 109 -23
rect 95 -37 99 -33
rect 114 -37 118 -9
rect 123 -21 127 -9
rect 123 -25 169 -21
rect 193 -25 197 -22
rect 165 -29 197 -25
rect 94 -41 99 -37
rect 108 -41 118 -37
rect 193 -35 197 -29
rect 201 -26 205 -22
rect 209 -26 213 -5
rect 240 -9 244 -5
rect 201 -30 213 -26
rect 225 -19 229 -16
rect 248 -19 252 -15
rect 278 -18 282 13
rect 225 -23 241 -19
rect 248 -23 265 -19
rect 278 -23 288 -18
rect 201 -35 205 -30
rect 95 -45 99 -41
rect 225 -45 229 -23
rect 248 -26 252 -23
rect 240 -32 244 -30
rect 105 -70 109 -49
rect 262 -54 266 -49
rect 147 -70 151 -54
rect 250 -58 266 -54
rect 240 -70 244 -67
rect 250 -70 254 -58
rect 262 -62 266 -58
rect 270 -53 274 -49
rect 278 -53 282 -23
rect 270 -57 282 -53
rect 270 -62 274 -57
rect -16 -74 254 -70
<< metal2 >>
rect 36 -19 40 3
rect 105 -19 109 3
rect 4 -37 8 -34
rect 73 -37 77 -34
rect 4 -41 21 -37
rect 73 -41 90 -37
rect 147 -50 151 0
rect 225 -12 229 35
rect 240 -63 244 -36
<< ntransistor >>
rect 152 6 154 10
rect 61 -2 63 6
rect -6 -20 -4 -12
rect 17 -16 19 -12
rect 86 -16 88 -12
rect 31 -49 35 -45
rect 267 3 269 9
rect 198 -3 200 3
rect 245 -30 247 -26
rect 198 -40 200 -34
rect 100 -49 104 -45
rect 267 -67 269 -61
<< ptransistor >>
rect -6 -2 -4 14
rect 152 20 154 28
rect 198 14 200 22
rect 267 20 269 28
rect 17 -2 19 6
rect 86 -2 88 6
rect 31 -34 35 -26
rect 61 -28 63 -12
rect 100 -34 104 -26
rect 198 -23 200 -15
rect 245 -16 247 -8
rect 267 -50 269 -42
<< polycontact >>
rect 265 35 269 39
rect 27 22 31 26
rect 148 13 152 17
rect 170 13 174 17
rect 13 -9 17 -5
rect 82 -9 86 -5
rect 35 -41 39 -37
rect 104 -41 108 -37
rect 196 -9 200 -5
rect 241 -23 245 -19
rect 265 -23 269 -19
rect 43 -67 47 -63
<< ndcontact >>
rect 147 6 151 10
rect 155 6 159 10
rect 56 -1 60 5
rect 64 -1 68 5
rect -11 -19 -7 -13
rect -3 -19 1 -13
rect 12 -16 16 -12
rect 20 -16 24 -12
rect 81 -16 85 -12
rect 89 -16 93 -12
rect 26 -49 30 -45
rect 36 -49 40 -45
rect 262 4 266 8
rect 270 4 274 8
rect 193 -2 197 2
rect 201 -2 205 2
rect 240 -30 244 -26
rect 248 -30 252 -26
rect 193 -39 197 -35
rect 201 -39 205 -35
rect 95 -49 99 -45
rect 105 -49 109 -45
rect 262 -66 266 -62
rect 270 -66 274 -62
<< pdcontact >>
rect -11 -1 -7 13
rect -3 -1 1 13
rect 147 21 151 27
rect 155 21 159 27
rect 193 15 197 21
rect 201 15 205 21
rect 262 21 266 27
rect 270 21 274 27
rect 12 -1 16 5
rect 20 -1 24 5
rect 81 -1 85 5
rect 89 -1 93 5
rect 26 -33 30 -27
rect 36 -33 40 -27
rect 56 -27 60 -13
rect 64 -27 68 -13
rect 95 -33 99 -27
rect 105 -33 109 -27
rect 240 -15 244 -9
rect 193 -22 197 -16
rect 248 -15 252 -9
rect 201 -22 205 -16
rect 262 -49 266 -43
rect 270 -49 274 -43
<< m2contact >>
rect 225 35 229 39
rect 36 3 40 7
rect 4 -34 8 -30
rect 36 -23 40 -19
rect 105 3 109 7
rect 147 0 151 4
rect 73 -34 77 -30
rect 21 -41 25 -37
rect 105 -23 109 -19
rect 90 -41 94 -37
rect 225 -16 229 -12
rect 240 -36 244 -32
rect 147 -54 151 -50
rect 240 -67 244 -63
<< labels >>
rlabel polycontact 27 22 31 26 0 clk
rlabel metal1 49 -9 56 -5 0 Qm
rlabel polycontact 43 -67 47 -63 0 not_clk
rlabel metal1 -13 -74 109 -70 0 gnd
rlabel metal1 -13 31 109 35 0 Vdd
rlabel metal1 -25 -10 -11 -5 0 D
rlabel metal1 132 -9 136 17 0 S
rlabel metal1 225 -45 229 -19 0 R
rlabel metal1 278 -23 288 -18 0 Q
<< end >>
