magic
tech scmos
timestamp 1672438776
<< polysilicon >>
rect -124 22 89 24
rect 93 22 240 24
rect -124 14 -122 22
rect 136 15 138 17
rect 79 6 81 8
rect -70 1 -68 3
rect 2 2 4 4
rect -124 -4 -122 -2
rect -124 -12 -122 -10
rect -124 -85 -122 -20
rect -93 -35 -91 -33
rect -93 -53 -91 -43
rect -70 -46 -68 -3
rect -56 -12 -54 -10
rect -56 -21 -54 -16
rect -56 -45 -54 -25
rect -25 -35 -23 -33
rect -70 -52 -68 -50
rect -25 -53 -23 -43
rect 2 -46 4 -2
rect 79 -12 81 -2
rect 13 -15 15 -12
rect 79 -18 81 -16
rect 2 -52 4 -50
rect -93 -59 -91 -57
rect -25 -59 -23 -57
rect 13 -59 15 -19
rect 93 -26 97 -24
rect 93 -45 97 -34
rect 136 -45 138 11
rect 238 6 240 22
rect 315 21 317 23
rect 315 0 317 13
rect 401 4 403 6
rect 238 -5 240 -2
rect 238 -12 240 -9
rect 315 -12 317 -4
rect 338 -6 360 -4
rect 150 -27 152 -25
rect 186 -28 188 -26
rect 93 -51 97 -49
rect 13 -64 15 -63
rect 136 -73 138 -49
rect 150 -54 152 -31
rect 150 -63 152 -58
rect 186 -76 188 -32
rect 199 -37 201 -36
rect 199 -44 201 -41
rect 199 -56 201 -48
rect 186 -83 188 -80
rect 238 -85 240 -28
rect 265 -46 267 -37
rect 255 -75 257 -65
rect 255 -82 257 -79
rect 265 -85 267 -50
rect 338 -61 340 -6
rect 358 -9 360 -6
rect 358 -16 360 -13
rect 401 -14 403 -4
rect 461 -13 463 -11
rect 401 -20 403 -18
rect 358 -23 360 -21
rect 415 -28 419 -26
rect 358 -33 360 -31
rect 461 -34 463 -21
rect 358 -47 360 -37
rect 415 -47 419 -36
rect 461 -46 463 -38
rect 358 -54 360 -51
rect 415 -53 419 -51
rect 358 -61 360 -59
rect 338 -73 340 -65
rect 358 -73 360 -69
rect 338 -75 360 -73
rect -124 -87 105 -85
rect 109 -87 240 -85
rect 265 -91 267 -89
<< ndiffusion >>
rect -76 -3 -75 1
rect -71 -3 -70 1
rect -68 -3 -67 1
rect -63 -3 -62 1
rect -4 -2 -3 2
rect 1 -2 2 2
rect 4 -2 5 2
rect 9 -2 10 2
rect -130 -13 -124 -12
rect -130 -19 -129 -13
rect -125 -19 -124 -13
rect -130 -20 -124 -19
rect -122 -13 -116 -12
rect -122 -19 -121 -13
rect -117 -19 -116 -13
rect -122 -20 -116 -19
rect -63 -16 -62 -12
rect -58 -16 -56 -12
rect -54 -16 -53 -12
rect -49 -16 -48 -12
rect 7 -19 8 -15
rect 12 -19 13 -15
rect 15 -19 16 -15
rect 20 -19 21 -15
rect 73 -16 74 -12
rect 78 -16 79 -12
rect 81 -16 82 -12
rect 86 -16 87 -12
rect -99 -57 -98 -53
rect -94 -57 -93 -53
rect -91 -57 -90 -53
rect -86 -57 -85 -53
rect -31 -57 -30 -53
rect -26 -57 -25 -53
rect -23 -57 -22 -53
rect -18 -57 -17 -53
rect 232 5 238 6
rect 232 -1 233 5
rect 237 -1 238 5
rect 232 -2 238 -1
rect 240 5 246 6
rect 240 -1 241 5
rect 245 -1 246 5
rect 240 -2 246 -1
rect 309 -4 310 0
rect 314 -4 315 0
rect 317 -4 318 0
rect 144 -31 145 -27
rect 149 -31 150 -27
rect 152 -31 153 -27
rect 157 -31 158 -27
rect 87 -49 88 -45
rect 92 -49 93 -45
rect 97 -49 98 -45
rect 102 -49 103 -45
rect 130 -49 131 -45
rect 135 -49 136 -45
rect 138 -49 139 -45
rect 143 -49 144 -45
rect 180 -32 181 -28
rect 185 -32 186 -28
rect 188 -32 189 -28
rect 193 -32 194 -28
rect 193 -48 194 -44
rect 198 -48 199 -44
rect 201 -48 202 -44
rect 206 -48 207 -44
rect 249 -79 250 -75
rect 254 -79 255 -75
rect 257 -79 258 -75
rect 262 -79 263 -75
rect 352 -13 353 -9
rect 357 -13 358 -9
rect 360 -13 361 -9
rect 365 -13 366 -9
rect 395 -18 396 -14
rect 400 -18 401 -14
rect 403 -18 404 -14
rect 408 -18 409 -14
rect 455 -38 456 -34
rect 460 -38 461 -34
rect 463 -38 464 -34
rect 352 -51 353 -47
rect 357 -51 358 -47
rect 360 -51 361 -47
rect 365 -51 366 -47
rect 409 -51 410 -47
rect 414 -51 415 -47
rect 419 -51 420 -47
rect 424 -51 425 -47
rect 259 -89 260 -85
rect 264 -89 265 -85
rect 267 -89 268 -85
rect 272 -89 273 -85
<< pdiffusion >>
rect -130 13 -124 14
rect -130 -1 -129 13
rect -125 -1 -124 13
rect -130 -2 -124 -1
rect -122 13 -116 14
rect -122 -1 -121 13
rect -117 -1 -116 13
rect 73 5 79 6
rect -122 -2 -116 -1
rect 73 -1 74 5
rect 78 -1 79 5
rect 73 -2 79 -1
rect 81 5 87 6
rect 81 -1 82 5
rect 86 -1 87 5
rect 81 -2 87 -1
rect -99 -36 -93 -35
rect -99 -42 -98 -36
rect -94 -42 -93 -36
rect -99 -43 -93 -42
rect -91 -36 -85 -35
rect -91 -42 -90 -36
rect -86 -42 -85 -36
rect -91 -43 -85 -42
rect -31 -36 -25 -35
rect -31 -42 -30 -36
rect -26 -42 -25 -36
rect -31 -43 -25 -42
rect -23 -36 -17 -35
rect -23 -42 -22 -36
rect -18 -42 -17 -36
rect -23 -43 -17 -42
rect 87 -27 93 -26
rect 87 -33 88 -27
rect 92 -33 93 -27
rect 87 -34 93 -33
rect 97 -27 103 -26
rect 97 -33 98 -27
rect 102 -33 103 -27
rect 97 -34 103 -33
rect 309 20 315 21
rect 309 14 310 20
rect 314 14 315 20
rect 309 13 315 14
rect 317 20 323 21
rect 317 14 318 20
rect 322 14 323 20
rect 317 13 323 14
rect 395 3 401 4
rect 395 -3 396 3
rect 400 -3 401 3
rect 395 -4 401 -3
rect 403 3 409 4
rect 403 -3 404 3
rect 408 -3 409 3
rect 403 -4 409 -3
rect 232 -13 238 -12
rect 232 -27 233 -13
rect 237 -27 238 -13
rect 232 -28 238 -27
rect 240 -13 246 -12
rect 240 -27 241 -13
rect 245 -27 246 -13
rect 240 -28 246 -27
rect 455 -14 461 -13
rect 455 -20 456 -14
rect 460 -20 461 -14
rect 455 -21 461 -20
rect 463 -14 469 -13
rect 463 -20 464 -14
rect 468 -20 469 -14
rect 463 -21 469 -20
rect 352 -24 358 -23
rect 352 -30 353 -24
rect 357 -30 358 -24
rect 352 -31 358 -30
rect 360 -24 366 -23
rect 360 -30 361 -24
rect 365 -30 366 -24
rect 360 -31 366 -30
rect 409 -29 415 -28
rect 409 -35 410 -29
rect 414 -35 415 -29
rect 409 -36 415 -35
rect 419 -29 425 -28
rect 419 -35 420 -29
rect 424 -35 425 -29
rect 419 -36 425 -35
rect 352 -62 358 -61
rect 352 -68 353 -62
rect 357 -68 358 -62
rect 352 -69 358 -68
rect 360 -62 366 -61
rect 360 -68 361 -62
rect 365 -68 366 -62
rect 360 -69 366 -68
<< metal1 >>
rect -131 31 460 35
rect -98 17 -94 31
rect -30 15 -26 31
rect -129 -5 -125 -1
rect -135 -9 -125 -5
rect -129 -13 -125 -9
rect 74 5 78 31
rect 98 7 102 31
rect 310 20 314 31
rect 118 11 135 15
rect 139 11 167 15
rect -121 -5 -117 -1
rect -110 -3 -75 1
rect -63 -3 -49 1
rect -110 -5 -106 -3
rect -121 -9 -106 -5
rect -53 -5 -49 -3
rect -10 -2 -3 2
rect 9 -2 26 2
rect 221 9 272 13
rect 318 9 322 14
rect -10 -5 -6 -2
rect -53 -9 -6 -5
rect 22 -5 26 -2
rect 82 -5 86 -1
rect 221 -5 226 9
rect 233 -5 237 -1
rect 22 -9 75 -5
rect 82 -9 237 -5
rect -121 -13 -117 -9
rect -114 -30 -110 -9
rect -53 -12 -49 -9
rect -78 -16 -62 -12
rect 22 -15 26 -9
rect 82 -12 86 -9
rect -78 -21 -74 -16
rect -7 -19 8 -15
rect 20 -19 26 -15
rect -105 -25 -57 -21
rect -105 -46 -101 -25
rect -98 -36 -94 -32
rect -90 -46 -86 -42
rect -107 -50 -97 -46
rect -90 -50 -71 -46
rect -90 -53 -86 -50
rect -98 -92 -94 -57
rect -80 -76 -76 -50
rect -64 -68 -60 -25
rect -30 -36 -26 -32
rect -22 -46 -18 -42
rect -7 -46 -3 -19
rect -43 -50 -29 -46
rect -22 -50 1 -46
rect 5 -50 26 -46
rect -42 -59 -38 -50
rect -22 -53 -18 -50
rect -30 -92 -26 -57
rect 33 -59 37 -20
rect 5 -63 12 -59
rect 16 -63 37 -59
rect 74 -92 78 -16
rect 98 -27 102 -23
rect 160 -24 178 -20
rect 160 -27 164 -24
rect 123 -31 145 -27
rect 157 -31 164 -27
rect 174 -28 178 -24
rect 204 -28 208 -9
rect 233 -13 237 -9
rect 241 -5 245 -1
rect 241 -9 257 -5
rect 241 -13 245 -9
rect 253 -24 257 -9
rect 268 -16 272 9
rect 299 5 311 9
rect 318 5 328 9
rect 318 0 322 5
rect 396 3 400 31
rect 420 5 424 31
rect 310 -9 314 -4
rect 404 -7 408 -3
rect 307 -13 314 -9
rect 353 -16 357 -13
rect 268 -20 357 -16
rect 353 -24 357 -20
rect 88 -37 92 -33
rect 123 -37 128 -31
rect 87 -41 92 -37
rect 101 -41 128 -37
rect 88 -45 92 -41
rect 123 -45 128 -41
rect 167 -45 171 -32
rect 123 -49 131 -45
rect 143 -49 171 -45
rect 174 -32 181 -28
rect 193 -32 208 -28
rect 253 -28 265 -24
rect 174 -44 178 -32
rect 195 -41 199 -37
rect 174 -48 194 -44
rect 198 -48 199 -44
rect 98 -92 102 -49
rect 110 -58 149 -54
rect 202 -59 206 -48
rect 173 -63 206 -59
rect 173 -69 177 -63
rect 214 -69 218 -59
rect 173 -73 218 -69
rect 221 -73 225 -41
rect 229 -43 246 -39
rect 229 -66 233 -43
rect 253 -54 257 -28
rect 361 -16 365 -13
rect 377 -11 397 -7
rect 404 -11 449 -7
rect 377 -16 381 -11
rect 404 -14 408 -11
rect 361 -20 381 -16
rect 361 -24 365 -20
rect 264 -43 274 -39
rect 270 -46 274 -43
rect 269 -50 274 -46
rect 295 -47 299 -30
rect 332 -33 349 -31
rect 332 -35 357 -33
rect 303 -47 307 -35
rect 345 -37 357 -35
rect 353 -54 357 -51
rect 253 -58 357 -54
rect 245 -61 249 -59
rect 245 -65 254 -61
rect 274 -65 337 -61
rect 353 -62 357 -58
rect 173 -76 177 -73
rect 221 -75 247 -73
rect 274 -75 278 -65
rect 361 -54 365 -51
rect 370 -54 374 -20
rect 361 -58 374 -54
rect 361 -62 365 -58
rect 295 -75 299 -74
rect 122 -80 185 -76
rect 221 -77 250 -75
rect 243 -79 250 -77
rect 262 -79 299 -75
rect 222 -85 226 -84
rect 274 -85 278 -79
rect 222 -89 260 -85
rect 272 -89 278 -85
rect 303 -92 307 -86
rect 396 -92 400 -18
rect 420 -29 424 -25
rect 410 -39 414 -35
rect 429 -39 433 -11
rect 445 -25 449 -11
rect 456 -14 460 31
rect 464 -25 468 -20
rect 445 -29 457 -25
rect 464 -29 477 -25
rect 464 -34 468 -29
rect 409 -43 414 -39
rect 423 -43 433 -39
rect 410 -47 414 -43
rect 420 -92 424 -51
rect 456 -92 460 -38
rect -128 -96 460 -92
<< metal2 >>
rect -98 -28 -94 13
rect -30 -28 -26 11
rect 33 11 114 15
rect 33 -16 37 11
rect 98 -19 102 3
rect 167 -13 171 11
rect 167 -17 217 -13
rect 167 -28 171 -17
rect -114 -37 -110 -34
rect 213 -37 217 -17
rect 269 -28 280 -24
rect -114 -41 83 -37
rect 111 -41 191 -37
rect 213 -41 221 -37
rect 277 -39 280 -28
rect 295 -26 299 5
rect 303 -31 307 -13
rect 328 -31 332 5
rect 420 -21 424 1
rect 30 -50 60 -46
rect 56 -54 60 -50
rect 56 -58 106 -54
rect -38 -63 1 -59
rect 116 -66 120 -41
rect 250 -43 260 -39
rect 277 -43 405 -39
rect 218 -59 245 -55
rect 31 -68 229 -66
rect -60 -70 229 -68
rect 295 -70 299 -51
rect -60 -72 34 -70
rect -76 -80 118 -76
rect 222 -80 226 -70
rect 303 -82 307 -51
<< ntransistor >>
rect -70 -3 -68 1
rect 2 -2 4 2
rect -124 -20 -122 -12
rect -56 -16 -54 -12
rect 13 -19 15 -15
rect 79 -16 81 -12
rect -93 -57 -91 -53
rect -25 -57 -23 -53
rect 238 -2 240 6
rect 315 -4 317 0
rect 150 -31 152 -27
rect 93 -49 97 -45
rect 136 -49 138 -45
rect 186 -32 188 -28
rect 199 -48 201 -44
rect 255 -79 257 -75
rect 358 -13 360 -9
rect 401 -18 403 -14
rect 461 -38 463 -34
rect 358 -51 360 -47
rect 415 -51 419 -47
rect 265 -89 267 -85
<< ptransistor >>
rect -124 -2 -122 14
rect 79 -2 81 6
rect -93 -43 -91 -35
rect -25 -43 -23 -35
rect 93 -34 97 -26
rect 315 13 317 21
rect 401 -4 403 4
rect 238 -28 240 -12
rect 461 -21 463 -13
rect 358 -31 360 -23
rect 415 -36 419 -28
rect 358 -69 360 -61
<< polycontact >>
rect 89 22 93 26
rect 135 11 139 15
rect -97 -50 -93 -46
rect -57 -25 -53 -21
rect -71 -50 -67 -46
rect -29 -50 -25 -46
rect 75 -9 79 -5
rect 1 -50 5 -46
rect 97 -41 101 -37
rect 311 5 315 9
rect 12 -63 16 -59
rect 149 -58 153 -54
rect 199 -41 203 -37
rect 185 -80 189 -76
rect 265 -50 269 -46
rect 254 -65 258 -61
rect 397 -11 401 -7
rect 357 -37 361 -33
rect 457 -29 461 -25
rect 419 -43 423 -39
rect 337 -65 341 -61
rect 105 -89 109 -85
<< ndcontact >>
rect -75 -3 -71 1
rect -67 -3 -63 1
rect -3 -2 1 2
rect 5 -2 9 2
rect -129 -19 -125 -13
rect -121 -19 -117 -13
rect -62 -16 -58 -12
rect -53 -16 -49 -12
rect 8 -19 12 -15
rect 16 -19 20 -15
rect 74 -16 78 -12
rect 82 -16 86 -12
rect -98 -57 -94 -53
rect -90 -57 -86 -53
rect -30 -57 -26 -53
rect -22 -57 -18 -53
rect 233 -1 237 5
rect 241 -1 245 5
rect 310 -4 314 0
rect 318 -4 322 0
rect 145 -31 149 -27
rect 153 -31 157 -27
rect 88 -49 92 -45
rect 98 -49 102 -45
rect 131 -49 135 -45
rect 139 -49 143 -45
rect 181 -32 185 -28
rect 189 -32 193 -28
rect 194 -48 198 -44
rect 202 -48 206 -44
rect 250 -79 254 -75
rect 258 -79 262 -75
rect 353 -13 357 -9
rect 361 -13 365 -9
rect 396 -18 400 -14
rect 404 -18 408 -14
rect 456 -38 460 -34
rect 464 -38 468 -34
rect 353 -51 357 -47
rect 361 -51 365 -47
rect 410 -51 414 -47
rect 420 -51 424 -47
rect 260 -89 264 -85
rect 268 -89 272 -85
<< pdcontact >>
rect -129 -1 -125 13
rect -121 -1 -117 13
rect 74 -1 78 5
rect 82 -1 86 5
rect -98 -42 -94 -36
rect -90 -42 -86 -36
rect -30 -42 -26 -36
rect -22 -42 -18 -36
rect 88 -33 92 -27
rect 98 -33 102 -27
rect 310 14 314 20
rect 318 14 322 20
rect 396 -3 400 3
rect 404 -3 408 3
rect 233 -27 237 -13
rect 241 -27 245 -13
rect 456 -20 460 -14
rect 464 -20 468 -14
rect 353 -30 357 -24
rect 361 -30 365 -24
rect 410 -35 414 -29
rect 420 -35 424 -29
rect 353 -68 357 -62
rect 361 -68 365 -62
<< m2contact >>
rect -98 13 -94 17
rect -30 11 -26 15
rect 114 11 118 15
rect 167 11 171 15
rect 98 3 102 7
rect -114 -34 -110 -30
rect -98 -32 -94 -28
rect -30 -32 -26 -28
rect 33 -20 37 -16
rect 26 -50 30 -46
rect -42 -63 -38 -59
rect -64 -72 -60 -68
rect -80 -80 -76 -76
rect 1 -63 5 -59
rect 98 -23 102 -19
rect 295 5 299 9
rect 328 5 332 9
rect 420 1 424 5
rect 303 -13 307 -9
rect 83 -41 87 -37
rect 167 -32 171 -28
rect 265 -28 269 -24
rect 191 -41 195 -37
rect 221 -41 225 -37
rect 106 -58 110 -54
rect 214 -59 218 -55
rect 246 -43 250 -39
rect 295 -30 299 -26
rect 260 -43 264 -39
rect 295 -51 299 -47
rect 303 -35 307 -31
rect 328 -35 332 -31
rect 303 -51 307 -47
rect 245 -59 249 -55
rect 229 -70 233 -66
rect 295 -74 299 -70
rect 118 -80 122 -76
rect 222 -84 226 -80
rect 303 -86 307 -82
rect 420 -25 424 -21
rect 405 -43 409 -39
<< labels >>
rlabel metal1 -135 -9 -129 -5 0 D
rlabel metal1 -107 -50 -99 -46 0 S
rlabel metal1 -114 -9 -106 -5 0 Dpass
rlabel metal1 -49 -9 -40 -5 0 or_1_out
rlabel metal1 -90 -50 -79 -46 0 not_S
rlabel metal1 207 -9 214 -5 0 Qm
rlabel metal1 245 -9 257 -5 0 Qpass
rlabel metal1 -43 -50 -31 -46 0 R
rlabel metal1 -22 -50 -10 -46 0 not_R
rlabel polycontact 105 -89 109 -85 0 not_clk
rlabel polycontact 89 22 93 26 0 clk
rlabel metal1 369 -20 381 -16 1 mux_out_1
rlabel metal1 433 -11 445 -7 0 Q
rlabel metal1 332 -35 349 -31 0 not_sel
rlabel metal1 263 -79 299 -75 0 sel
rlabel metal1 468 -29 477 -25 0 Qbar
rlabel metal1 -131 31 460 35 0 Vdd
rlabel metal1 -128 -96 460 -92 0 gnd
<< end >>
